package sharedpkg ;
parameter FIFO_WIDTH = 16;
parameter FIFO_DEPTH = 8;
int error_count = 0  ;
int correct_count = 0; 
    
endpackage